`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:46:45 10/08/2022 
// Design Name: 
// Module Name:    dec_gray532_bh 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

// AYUSH GUPTA
// Gray Code to Unsigned Thermometer Code Decoder

// NOTE : 5-bit Input Gray Code
// 	  : 32 bits Output Thermometer code with MSB as Unsigned Bit

module dec_gray532_bh
(
	input      [4:0]  I,
	output reg [31:0] O
);

always @(I)
begin

	case (I)
		5'b00000 : O = 32'b00000000000000000000000000000000;
		5'b00001 : O = 32'b00000000000000000000000000000001;
		5'b00011 : O = 32'b00000000000000000000000000000011;
		5'b00010 : O = 32'b00000000000000000000000000000111;
		5'b00110 : O = 32'b00000000000000000000000000001111;
		5'b00111 : O = 32'b00000000000000000000000000011111;
		5'b00101 : O = 32'b00000000000000000000000000111111;
		5'b00100 : O = 32'b00000000000000000000000001111111;
		5'b01100 : O = 32'b00000000000000000000000011111111;
		5'b01101 : O = 32'b00000000000000000000000111111111;
		5'b01111 : O = 32'b00000000000000000000001111111111;
		5'b01110 : O = 32'b00000000000000000000011111111111;
		5'b01010 : O = 32'b00000000000000000000111111111111;
		5'b01011 : O = 32'b00000000000000000001111111111111;
		5'b01001 : O = 32'b00000000000000000011111111111111;
		5'b01000 : O = 32'b00000000000000000111111111111111;
		5'b11000 : O = 32'b00000000000000001111111111111111;
		5'b11001 : O = 32'b00000000000000011111111111111111;
		5'b11011 : O = 32'b00000000000000111111111111111111;
		5'b11010 : O = 32'b00000000000001111111111111111111;
		5'b11110 : O = 32'b00000000000011111111111111111111;
		5'b11111 : O = 32'b00000000000111111111111111111111;
		5'b11101 : O = 32'b00000000001111111111111111111111;
		5'b11100 : O = 32'b00000000011111111111111111111111;
		5'b10100 : O = 32'b00000000111111111111111111111111;
		5'b10101 : O = 32'b00000001111111111111111111111111;
		5'b10111 : O = 32'b00000011111111111111111111111111;
		5'b10110 : O = 32'b00000111111111111111111111111111;
		5'b10010 : O = 32'b00001111111111111111111111111111;
		5'b10011 : O = 32'b00011111111111111111111111111111;
		5'b10001 : O = 32'b00111111111111111111111111111111;
		5'b10000 : O = 32'b01111111111111111111111111111111;
	   default  : O = "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";
	 endcase
	 
end
endmodule
